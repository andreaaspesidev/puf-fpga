`timescale 1ns / 1ps

module tb_CompFreq;

  reg clk = 0;
  
  reg [7:0] challenge;
  reg increment = 0;
  reg reset = 0;
  reg [10:0] nextT;
  reg done;
  //reg [7:0] conf;
  reg [10:0] count;

  //reg [7:0] challenge14_indices [0:119] = {8'd1, 8'd2, 8'd3, 8'd4, 8'd5, 8'd6, 8'd7, 8'd8, 8'd9, 8'd10, 8'd11, 8'd12, 8'd13, 8'd14, 8'd15, 8'd239, 8'd18, 8'd19, 8'd20, 8'd21, 8'd22, 8'd23, 8'd24, 8'd25, 8'd26, 8'd27, 8'd28, 8'd29, 8'd30, 8'd31, 8'd222, 8'd223, 8'd35, 8'd36, 8'd37, 8'd38, 8'd39, 8'd40, 8'd41, 8'd42, 8'd43, 8'd44, 8'd45, 8'd46, 8'd47, 8'd205, 8'd206, 8'd207, 8'd52, 8'd53, 8'd54, 8'd55, 8'd56, 8'd57, 8'd58, 8'd59, 8'd60, 8'd61, 8'd62, 8'd63, 8'd188, 8'd189, 8'd190, 8'd191, 8'd69, 8'd70, 8'd71, 8'd72, 8'd73, 8'd74, 8'd75, 8'd76, 8'd77, 8'd78, 8'd79, 8'd171, 8'd172, 8'd173, 8'd174, 8'd175, 8'd86, 8'd87, 8'd88, 8'd89, 8'd90, 8'd91, 8'd92, 8'd93, 8'd94, 8'd95, 8'd154, 8'd155, 8'd156, 8'd157, 8'd158, 8'd159, 8'd103, 8'd104, 8'd105, 8'd106, 8'd107, 8'd108, 8'd109, 8'd110, 8'd111, 8'd137, 8'd138, 8'd139, 8'd140, 8'd141, 8'd142, 8'd143, 8'd120, 8'd121, 8'd122, 8'd123, 8'd124, 8'd125, 8'd126, 8'd127};
  reg [10:0] challenge14_freqs [0:159] = {11'd0, 11'd128, 11'd256, 11'd384, 11'd512, 11'd640, 11'd768, 11'd896, 11'd1024, 11'd1152, 11'd1, 11'd129, 11'd257, 11'd385, 11'd513, 11'd641, 11'd769, 11'd897, 11'd1025, 11'd1153, 11'd2, 11'd130, 11'd258, 11'd386, 11'd514, 11'd642, 11'd770, 11'd898, 11'd1026, 11'd1154, 11'd3, 11'd131, 11'd259, 11'd387, 11'd515, 11'd643, 11'd771, 11'd899, 11'd1027, 11'd1155, 11'd4, 11'd132, 11'd260, 11'd388, 11'd516, 11'd644, 11'd772, 11'd900, 11'd1028, 11'd1156, 11'd5, 11'd133, 11'd261, 11'd389, 11'd517, 11'd645, 11'd773, 11'd901, 11'd1029, 11'd1157, 11'd6, 11'd134, 11'd262, 11'd390, 11'd518, 11'd646, 11'd774, 11'd902, 11'd1030, 11'd1158, 11'd7, 11'd135, 11'd263, 11'd391, 11'd519, 11'd647, 11'd775, 11'd903, 11'd1031, 11'd1159, 11'd120, 11'd248, 11'd376, 11'd504, 11'd632, 11'd760, 11'd888, 11'd1016, 11'd1144, 11'd1272, 11'd121, 11'd249, 11'd377, 11'd505, 11'd633, 11'd761, 11'd889, 11'd1017, 11'd1145, 11'd1273, 11'd122, 11'd250, 11'd378, 11'd506, 11'd634, 11'd762, 11'd890, 11'd1018, 11'd1146, 11'd1274, 11'd123, 11'd251, 11'd379, 11'd507, 11'd635, 11'd763, 11'd891, 11'd1019, 11'd1147, 11'd1275, 11'd124, 11'd252, 11'd380, 11'd508, 11'd636, 11'd764, 11'd892, 11'd1020, 11'd1148, 11'd1276, 11'd125, 11'd253, 11'd381, 11'd509, 11'd637, 11'd765, 11'd893, 11'd1021, 11'd1149, 11'd1277, 11'd126, 11'd254, 11'd382, 11'd510, 11'd638, 11'd766, 11'd894, 11'd1022, 11'd1150, 11'd1278, 11'd127, 11'd255, 11'd383, 11'd511, 11'd639, 11'd767, 11'd895, 11'd1023, 11'd1151, 11'd1279};
  reg [10:0] challenge58_freqs [0:159] = {11'd24, 11'd152, 11'd280, 11'd408, 11'd536, 11'd664, 11'd792, 11'd920, 11'd1048, 11'd1176, 11'd25, 11'd153, 11'd281, 11'd409, 11'd537, 11'd665, 11'd793, 11'd921, 11'd1049, 11'd1177, 11'd26, 11'd154, 11'd282, 11'd410, 11'd538, 11'd666, 11'd794, 11'd922, 11'd1050, 11'd1178, 11'd27, 11'd155, 11'd283, 11'd411, 11'd539, 11'd667, 11'd795, 11'd923, 11'd1051, 11'd1179, 11'd28, 11'd156, 11'd284, 11'd412, 11'd540, 11'd668, 11'd796, 11'd924, 11'd1052, 11'd1180, 11'd29, 11'd157, 11'd285, 11'd413, 11'd541, 11'd669, 11'd797, 11'd925, 11'd1053, 11'd1181, 11'd30, 11'd158, 11'd286, 11'd414, 11'd542, 11'd670, 11'd798, 11'd926, 11'd1054, 11'd1182, 11'd31, 11'd159, 11'd287, 11'd415, 11'd543, 11'd671, 11'd799, 11'd927, 11'd1055, 11'd1183, 11'd112, 11'd240, 11'd368, 11'd496, 11'd624, 11'd752, 11'd880, 11'd1008, 11'd1136, 11'd1264, 11'd113, 11'd241, 11'd369, 11'd497, 11'd625, 11'd753, 11'd881, 11'd1009, 11'd1137, 11'd1265, 11'd114, 11'd242, 11'd370, 11'd498, 11'd626, 11'd754, 11'd882, 11'd1010, 11'd1138, 11'd1266, 11'd115, 11'd243, 11'd371, 11'd499, 11'd627, 11'd755, 11'd883, 11'd1011, 11'd1139, 11'd1267, 11'd116, 11'd244, 11'd372, 11'd500, 11'd628, 11'd756, 11'd884, 11'd1012, 11'd1140, 11'd1268, 11'd117, 11'd245, 11'd373, 11'd501, 11'd629, 11'd757, 11'd885, 11'd1013, 11'd1141, 11'd1269, 11'd118, 11'd246, 11'd374, 11'd502, 11'd630, 11'd758, 11'd886, 11'd1014, 11'd1142, 11'd1270, 11'd119, 11'd247, 11'd375, 11'd503, 11'd631, 11'd759, 11'd887, 11'd1015, 11'd1143, 11'd1271};  
  reg [10:0] challenge61_freqs [0:159] = {11'd88, 11'd216, 11'd344, 11'd472, 11'd600, 11'd728, 11'd856, 11'd984, 11'd1112, 11'd1240, 11'd89, 11'd217, 11'd345, 11'd473, 11'd601, 11'd729, 11'd857, 11'd985, 11'd1113, 11'd1241, 11'd90, 11'd218, 11'd346, 11'd474, 11'd602, 11'd730, 11'd858, 11'd986, 11'd1114, 11'd1242, 11'd91, 11'd219, 11'd347, 11'd475, 11'd603, 11'd731, 11'd859, 11'd987, 11'd1115, 11'd1243, 11'd92, 11'd220, 11'd348, 11'd476, 11'd604, 11'd732, 11'd860, 11'd988, 11'd1116, 11'd1244, 11'd93, 11'd221, 11'd349, 11'd477, 11'd605, 11'd733, 11'd861, 11'd989, 11'd1117, 11'd1245, 11'd94, 11'd222, 11'd350, 11'd478, 11'd606, 11'd734, 11'd862, 11'd990, 11'd1118, 11'd1246, 11'd95, 11'd223, 11'd351, 11'd479, 11'd607, 11'd735, 11'd863, 11'd991, 11'd1119, 11'd1247, 11'd104, 11'd232, 11'd360, 11'd488, 11'd616, 11'd744, 11'd872, 11'd1000, 11'd1128, 11'd1256, 11'd105, 11'd233, 11'd361, 11'd489, 11'd617, 11'd745, 11'd873, 11'd1001, 11'd1129, 11'd1257, 11'd106, 11'd234, 11'd362, 11'd490, 11'd618, 11'd746, 11'd874, 11'd1002, 11'd1130, 11'd1258, 11'd107, 11'd235, 11'd363, 11'd491, 11'd619, 11'd747, 11'd875, 11'd1003, 11'd1131, 11'd1259, 11'd108, 11'd236, 11'd364, 11'd492, 11'd620, 11'd748, 11'd876, 11'd1004, 11'd1132, 11'd1260, 11'd109, 11'd237, 11'd365, 11'd493, 11'd621, 11'd749, 11'd877, 11'd1005, 11'd1133, 11'd1261, 11'd110, 11'd238, 11'd366, 11'd494, 11'd622, 11'd750, 11'd878, 11'd1006, 11'd1134, 11'd1262, 11'd111, 11'd239, 11'd367, 11'd495, 11'd623, 11'd751, 11'd879, 11'd1007, 11'd1135, 11'd1263};

  comp_freq_cnt comp_freq_inst (
    .clk(clk),
    .challenge_in(challenge),
    .increment(increment),
    .reset(reset),
    .next_TERO(nextT),
    .done(done)
  );

  //assign conf = {comp_freq_inst.i, comp_freq_inst.j};

  initial begin
    begin
        clk <= 0;
        reset = 1;
        count = 0;
        increment = 0;
        // Inspect i,j are correctly generated
        //for (challenge = 0; challenge < 120; challenge = challenge + 1) begin
        //  @(posedge(clk));
        //  assert (conf == challenge_indices[challenge]);
        //end
        
        // Inspect frequencies outputs for challenge 14
        challenge = 14;
        reset = 1;
        repeat(20) @(posedge(clk));
        reset = 0;
        count = 0;
        @(posedge(clk));
        
        repeat (170) begin
          if (nextT != challenge14_freqs[count]) begin
            $display("[%d] %d %d\n", count, challenge14_freqs[count], nextT);
            $finish;
          end
          increment = 1;
          @(posedge(clk));
          increment = 0;
          @(posedge(clk));
          count = count + 1;
        end
        
        // Test second round, challenge 14
        reset = 1;
        repeat(20) @(posedge(clk));
        reset = 0;
        count = 0;
        @(posedge(clk));
        
        repeat (170) begin
          if (nextT != challenge14_freqs[count]) begin
            $display("[%d] %d %d\n", count, challenge14_freqs[count], nextT);
            $finish;
          end
          increment = 1;
          @(posedge(clk));
          increment = 0;
          @(posedge(clk));
          count = count + 1;
        end
        
        // Test challenge 58
        challenge = 58;
        reset = 1;
        repeat(20) @(posedge(clk));
        reset = 0;
        count = 0;
        @(posedge(clk));
        
        repeat (170) begin
          if (nextT != challenge58_freqs[count]) begin
            $display("[%d] %d %d\n", count, challenge58_freqs[count], nextT);
            $finish;
          end
          increment = 1;
          @(posedge(clk));
          increment = 0;
          @(posedge(clk));
          count = count + 1;
        end
        
        // Test challenge 61
        challenge = 61;
        reset = 1;
        repeat(20) @(posedge(clk));
        reset = 0;
        count = 0;
        @(posedge(clk));
        
        repeat (170) begin
          if (nextT != challenge61_freqs[count]) begin
            $display("[%d] %d %d\n", count, challenge61_freqs[count], nextT);
            $finish;
          end
          increment = 1;
          @(posedge(clk));
          increment = 0;
          @(posedge(clk));
          count = count + 1;
        end
        

      $finish; //end the simulation
    end
  end

  always
    #5  clk =~ clk ;

endmodule
